Starta från hårddisk Startalternativ Avbryt Ändra startdisk Fortsätt Katalog
 Uppdatera drivrutin Ha disketten för drivrutinsuppdatering redo. 

Det verkar som systemet startade från den andra sidan på dvd:n.
Om så är fallet, vänd på dvd:n och försök igen. Det här är en dvd med två sidor. Du har startat från den andra sidan.

Vänd på dvd:n och fortsätt sedan. Du är nästan klar... I/O-fel Du är på väg att lämna den grafiska startmenyn och
starta textlägesgränssnittet. Hej då FTP-installation Hårddisk Hårddiskinstallation Diskenhet (avsök alla diskar om tom)
 Hjälp HTTP-installation Starthanterare Sätt i startdisk %u. Det här är startdisk %u.
Sätt i startdisk %u. Det här är inte en Suse Linux 9.1-startdisk.
Sätt i startdisk %u. Installation Laddar Linux-kärna


 Startar... Laddar memtest86


 Manuell installation Minnestest NFS-installation Installation - ACPI inaktiverat OK Lösenord
 Lösenord Vill du stänga av systemet nu? Stäng av Starta om Räddningssystem Installation - Säkra inställningar Linux - Säkra inställningar Server
 SMB- (Windows-utdelning) installation Användare (anonym inloggning om tom)
 Användare (använder \"guest\" om tom)
 